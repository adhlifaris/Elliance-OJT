

///////////
//Central Control Fabric
//////////

//=====//
// System Control
//=====//

//=====//
//Clock Domain Manager
//=====//

//=====//
//Power Mode Controller 
//=====//
//////////////
// Config and Control Subsystem
//////////////

//////////
// Compute Cluster Array
/////////

////////
//Memory Subsystem
///////

////////
//Data Movement Engine
////////

///////
//Power Management Subsystem
//////

//////
//External Imterface
/////

////
//Monitoring and Telemetry
///

